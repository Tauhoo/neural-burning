module mult_matrix_prep(input_stream, output_stream, clk);

endmodule
