// data_path.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module data_path (
		input  wire        clk_clk,                                                      //                                               clk.clk
		input  wire        code_storage_code_control_interface_active,                   //               code_storage_code_control_interface.active
		input  wire        code_storage_code_control_interface_reset,                    //                                                  .reset
		input  wire [11:0] code_storage_write_interface_write_data,                      //                      code_storage_write_interface.write_data
		input  wire        code_storage_write_interface_is_write,                        //                                                  .is_write
		input  wire [31:0] code_storage_write_interface_write_line,                      //                                                  .write_line
		output wire [31:0] fetch_to_decode_register_code_index_out_interface_code_index, // fetch_to_decode_register_code_index_out_interface.code_index
		output wire        parse_clock_source_clk,                                       //                                parse_clock_source.clk
		output wire [3:0]  parse_op_interface_op,                                        //                                parse_op_interface.op
		output wire [3:0]  parse_parameter_type_interface_act_type,                      //                    parse_parameter_type_interface.act_type
		output wire [3:0]  parse_parameter_type_interface_dense_type,                    //                                                  .dense_type
		output wire [7:0]  parse_parameter_type_interface_cost_type,                     //                                                  .cost_type
		input  wire        reset_reset_n                                                 //                                             reset.reset_n
	);

	wire         fetch_to_decode_register_clock_source_clk;        // fetch_to_decode_register:clk_out -> parse:clk
	wire         code_storage_clock_source_clk;                    // code_storage:clk_out -> fetch_to_decode_register:clk
	wire  [11:0] code_storage_code_interface_code;                 // code_storage:code -> fetch_to_decode_register:code
	wire  [31:0] code_storage_code_interface_code_index;           // code_storage:code_index -> fetch_to_decode_register:code_index
	wire  [11:0] fetch_to_decode_register_code_out_interface_code; // fetch_to_decode_register:code_out -> parse:code

	code_storage #(
		.code_size     (12),
		.max_code_line (100)
	) code_storage (
		.clk        (clk_clk),                                    //                  clock.clk
		.code       (code_storage_code_interface_code),           //         code_interface.code
		.code_index (code_storage_code_interface_code_index),     //                       .code_index
		.active     (code_storage_code_control_interface_active), // code_control_interface.active
		.reset      (code_storage_code_control_interface_reset),  //                       .reset
		.write_data (code_storage_write_interface_write_data),    //        write_interface.write_data
		.is_write   (code_storage_write_interface_is_write),      //                       .is_write
		.write_line (code_storage_write_interface_write_line),    //                       .write_line
		.clk_out    (code_storage_clock_source_clk)               //           clock_source.clk
	);

	fetch_decode_reg #(
		.code_size (12)
	) fetch_to_decode_register (
		.clk            (code_storage_clock_source_clk),                                //                    clock.clk
		.code           (code_storage_code_interface_code),                             //           code_interface.code
		.code_index     (code_storage_code_interface_code_index),                       //                         .code_index
		.code_out       (fetch_to_decode_register_code_out_interface_code),             //       code_out_interface.code
		.code_index_out (fetch_to_decode_register_code_index_out_interface_code_index), // code_index_out_interface.code_index
		.clk_out        (fetch_to_decode_register_clock_source_clk)                     //             clock_source.clk
	);

	parse #(
		.op_size      (4),
		.param_a_size (4),
		.param_b_size (4)
	) parse (
		.code       (fetch_to_decode_register_code_out_interface_code), //           code_interface.code
		.act_type   (parse_parameter_type_interface_act_type),          // parameter_type_interface.act_type
		.dense_type (parse_parameter_type_interface_dense_type),        //                         .dense_type
		.cost_type  (parse_parameter_type_interface_cost_type),         //                         .cost_type
		.op         (parse_op_interface_op),                            //             op_interface.op
		.clk        (fetch_to_decode_register_clock_source_clk),        //                    clock.clk
		.clk_out    (parse_clock_source_clk)                            //             clock_source.clk
	);

endmodule
