module register_delay();
endmodule
